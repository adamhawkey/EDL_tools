<ColorDecisionList xmnls="urn:ASC:CDL:v1.01">
    <ColorDecision>
        <ColorCorrection>
            <SOPNode>
                <Slope>0.9330 0.9330 0.9244</Slope>
                <Offset>0.0671 0.0670 0.0755</Offset>
                <Power>1.0000 1.0000 1.0000</Power>
            </SOPNode>
            <SatNode>
                <Saturation>1.0000</Saturation>
            </SatNode>
        </ColorCorrection>
    </ColorDecision>
</ColorDecisionList>
