<?xml version="1.0" encoding="UTF-8"?>
<ViewingDescription>written with CDL_extract_0.2 by Adam Hawkey</ViewingDescription>
<ColorDecisionList xmnls="urn:ASC:CDL:v1.01">
    <ColorDecision>
        <ColorCorrection>
            <SOPNode>
                <Slope>0.927994 0.934545 1.043792</Slope>
                <Offset>0.065299 0.0554 -0.049585</Offset>
                <Power>1.055597 1.094934 0.967334</Power>
            </SOPNode>
            <SatNode>
                <Saturation>1.246499</Saturation>
            </SatNode>
        </ColorCorrection>
    </ColorDecision>
</ColorDecisionList>
